`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Create by Engineer: yaxingshi
// Create Date: 2023-03-24 15:11:30
// Last Modified by:   yaxingshi
// Last Modified time: 2023-03-24 15:32:41
// Design Name: 
// Module Name: line_delay_cal
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module line_delay_cal (
	input clk,    // Clock
	input rst,  // Asynchronous reset active low
	input 
	
);

endmodule : line_delay_cal